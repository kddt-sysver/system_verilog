module twd1_64 (
    input logic [8:0] rom_address_in, // 0에서 511까지의 단일 인덱스 입력
    output logic signed [8:0] twf_re_out,
    output logic signed [8:0] twf_im_out
);
    parameter int DATA_WIDTH = 9;  // Total bits for <2.7> (signed [8:0])
    parameter int ROM_DEPTH = 64;  // 8 * 8
    logic signed [DATA_WIDTH-1:0] twf_m1_re_rom[ROM_DEPTH-1:0];
    logic signed [DATA_WIDTH-1:0] twf_m1_im_rom[ROM_DEPTH-1:0];
    assign twf_re_out = twf_m1_re_rom[rom_address_in];
    assign twf_im_out = twf_m1_im_rom[rom_address_in];
    assign twf_m1_re_rom[0] = 128;
    assign twf_m1_im_rom[0] = 0;
    assign twf_m1_re_rom[1] = 128;
    assign twf_m1_im_rom[1] = 0;
    assign twf_m1_re_rom[2] = 128;
    assign twf_m1_im_rom[2] = 0;
    assign twf_m1_re_rom[3] = 128;
    assign twf_m1_im_rom[3] = 0;
    assign twf_m1_re_rom[4] = 128;
    assign twf_m1_im_rom[4] = 0;
    assign twf_m1_re_rom[5] = 128;
    assign twf_m1_im_rom[5] = 0;
    assign twf_m1_re_rom[6] = 128;
    assign twf_m1_im_rom[6] = 0;
    assign twf_m1_re_rom[7] = 128;
    assign twf_m1_im_rom[7] = 0;
    assign twf_m1_re_rom[8] = 128;
    assign twf_m1_im_rom[8] = 0;
    assign twf_m1_re_rom[9] = 118;
    assign twf_m1_im_rom[9] = -49;
    assign twf_m1_re_rom[10] = 91;
    assign twf_m1_im_rom[10] = -91;
    assign twf_m1_re_rom[11] = 49;
    assign twf_m1_im_rom[11] = -118;
    assign twf_m1_re_rom[12] = 0;
    assign twf_m1_im_rom[12] = -128;
    assign twf_m1_re_rom[13] = -49;
    assign twf_m1_im_rom[13] = -118;
    assign twf_m1_re_rom[14] = -91;
    assign twf_m1_im_rom[14] = -91;
    assign twf_m1_re_rom[15] = -118;
    assign twf_m1_im_rom[15] = -49;
    assign twf_m1_re_rom[16] = 128;
    assign twf_m1_im_rom[16] = 0;
    assign twf_m1_re_rom[17] = 126;
    assign twf_m1_im_rom[17] = -25;
    assign twf_m1_re_rom[18] = 118;
    assign twf_m1_im_rom[18] = -49;
    assign twf_m1_re_rom[19] = 106;
    assign twf_m1_im_rom[19] = -71;
    assign twf_m1_re_rom[20] = 91;
    assign twf_m1_im_rom[20] = -91;
    assign twf_m1_re_rom[21] = 71;
    assign twf_m1_im_rom[21] = -106;
    assign twf_m1_re_rom[22] = 49;
    assign twf_m1_im_rom[22] = -118;
    assign twf_m1_re_rom[23] = 25;
    assign twf_m1_im_rom[23] = -126;
    assign twf_m1_re_rom[24] = 128;
    assign twf_m1_im_rom[24] = 0;
    assign twf_m1_re_rom[25] = 106;
    assign twf_m1_im_rom[25] = -71;
    assign twf_m1_re_rom[26] = 49;
    assign twf_m1_im_rom[26] = -118;
    assign twf_m1_re_rom[27] = -25;
    assign twf_m1_im_rom[27] = -126;
    assign twf_m1_re_rom[28] = -91;
    assign twf_m1_im_rom[28] = -91;
    assign twf_m1_re_rom[29] = -126;
    assign twf_m1_im_rom[29] = -25;
    assign twf_m1_re_rom[30] = -118;
    assign twf_m1_im_rom[30] = 49;
    assign twf_m1_re_rom[31] = -71;
    assign twf_m1_im_rom[31] = 106;
    assign twf_m1_re_rom[32] = 128;
    assign twf_m1_im_rom[32] = 0;
    assign twf_m1_re_rom[33] = 127;
    assign twf_m1_im_rom[33] = -13;
    assign twf_m1_re_rom[34] = 126;
    assign twf_m1_im_rom[34] = -25;
    assign twf_m1_re_rom[35] = 122;
    assign twf_m1_im_rom[35] = -37;
    assign twf_m1_re_rom[36] = 118;
    assign twf_m1_im_rom[36] = -49;
    assign twf_m1_re_rom[37] = 113;
    assign twf_m1_im_rom[37] = -60;
    assign twf_m1_re_rom[38] = 106;
    assign twf_m1_im_rom[38] = -71;
    assign twf_m1_re_rom[39] = 99;
    assign twf_m1_im_rom[39] = -81;
    assign twf_m1_re_rom[40] = 128;
    assign twf_m1_im_rom[40] = 0;
    assign twf_m1_re_rom[41] = 113;
    assign twf_m1_im_rom[41] = -60;
    assign twf_m1_re_rom[42] = 71;
    assign twf_m1_im_rom[42] = -106;
    assign twf_m1_re_rom[43] = 13;
    assign twf_m1_im_rom[43] = -127;
    assign twf_m1_re_rom[44] = -49;
    assign twf_m1_im_rom[44] = -118;
    assign twf_m1_re_rom[45] = -99;
    assign twf_m1_im_rom[45] = -81;
    assign twf_m1_re_rom[46] = -126;
    assign twf_m1_im_rom[46] = -25;
    assign twf_m1_re_rom[47] = -122;
    assign twf_m1_im_rom[47] = 37;
    assign twf_m1_re_rom[48] = 128;
    assign twf_m1_im_rom[48] = 0;
    assign twf_m1_re_rom[49] = 122;
    assign twf_m1_im_rom[49] = -37;
    assign twf_m1_re_rom[50] = 106;
    assign twf_m1_im_rom[50] = -71;
    assign twf_m1_re_rom[51] = 81;
    assign twf_m1_im_rom[51] = -99;
    assign twf_m1_re_rom[52] = 49;
    assign twf_m1_im_rom[52] = -118;
    assign twf_m1_re_rom[53] = 13;
    assign twf_m1_im_rom[53] = -127;
    assign twf_m1_re_rom[54] = -25;
    assign twf_m1_im_rom[54] = -126;
    assign twf_m1_re_rom[55] = -60;
    assign twf_m1_im_rom[55] = -113;
    assign twf_m1_re_rom[56] = 128;
    assign twf_m1_im_rom[56] = 0;
    assign twf_m1_re_rom[57] = 99;
    assign twf_m1_im_rom[57] = -81;
    assign twf_m1_re_rom[58] = 25;
    assign twf_m1_im_rom[58] = -126;
    assign twf_m1_re_rom[59] = -60;
    assign twf_m1_im_rom[59] = -113;
    assign twf_m1_re_rom[60] = -118;
    assign twf_m1_im_rom[60] = -49;
    assign twf_m1_re_rom[61] = -122;
    assign twf_m1_im_rom[61] = 37;
    assign twf_m1_re_rom[62] = -71;
    assign twf_m1_im_rom[62] = 106;
    assign twf_m1_re_rom[63] = 13;
    assign twf_m1_im_rom[63] = 127;

endmodule
