module twd0_512 (
    input logic [8:0] rom_address_in, // 0에서 511까지의 단일 인덱스 입력
    output logic signed [8:0] twf_re_out,
    output logic signed [8:0] twf_im_out
);

    // --- Parameters and Constants ---
    parameter int DATA_WIDTH = 9;  // Total bits for <2.7> (signed [8:0])
    parameter int ROM_DEPTH = 512;  // 8 * 64

    // ROM arrays for real and imaginary parts
    // 이 배열들은 툴에 의해 BRAM (Block RAM)으로 합성될 수 있습니다.
    logic signed [DATA_WIDTH-1:0] twf_m0_re_rom[ROM_DEPTH-1:0];
    logic signed [DATA_WIDTH-1:0] twf_m0_im_rom[ROM_DEPTH-1:0];

    assign twf_re_out = twf_m0_re_rom[rom_address_in];
    assign twf_im_out = twf_m0_im_rom[rom_address_in];
    assign twf_m0_re_rom[0] = 128;
    assign twf_m0_im_rom[0] = 0;
    assign twf_m0_re_rom[1] = 128;
    assign twf_m0_im_rom[1] = 0;
    assign twf_m0_re_rom[2] = 128;
    assign twf_m0_im_rom[2] = 0;
    assign twf_m0_re_rom[3] = 128;
    assign twf_m0_im_rom[3] = 0;
    assign twf_m0_re_rom[4] = 128;
    assign twf_m0_im_rom[4] = 0;
    assign twf_m0_re_rom[5] = 128;
    assign twf_m0_im_rom[5] = 0;
    assign twf_m0_re_rom[6] = 128;
    assign twf_m0_im_rom[6] = 0;
    assign twf_m0_re_rom[7] = 128;
    assign twf_m0_im_rom[7] = 0;
    assign twf_m0_re_rom[8] = 128;
    assign twf_m0_im_rom[8] = 0;
    assign twf_m0_re_rom[9] = 128;
    assign twf_m0_im_rom[9] = 0;
    assign twf_m0_re_rom[10] = 128;
    assign twf_m0_im_rom[10] = 0;
    assign twf_m0_re_rom[11] = 128;
    assign twf_m0_im_rom[11] = 0;
    assign twf_m0_re_rom[12] = 128;
    assign twf_m0_im_rom[12] = 0;
    assign twf_m0_re_rom[13] = 128;
    assign twf_m0_im_rom[13] = 0;
    assign twf_m0_re_rom[14] = 128;
    assign twf_m0_im_rom[14] = 0;
    assign twf_m0_re_rom[15] = 128;
    assign twf_m0_im_rom[15] = 0;
    assign twf_m0_re_rom[16] = 128;
    assign twf_m0_im_rom[16] = 0;
    assign twf_m0_re_rom[17] = 128;
    assign twf_m0_im_rom[17] = 0;
    assign twf_m0_re_rom[18] = 128;
    assign twf_m0_im_rom[18] = 0;
    assign twf_m0_re_rom[19] = 128;
    assign twf_m0_im_rom[19] = 0;
    assign twf_m0_re_rom[20] = 128;
    assign twf_m0_im_rom[20] = 0;
    assign twf_m0_re_rom[21] = 128;
    assign twf_m0_im_rom[21] = 0;
    assign twf_m0_re_rom[22] = 128;
    assign twf_m0_im_rom[22] = 0;
    assign twf_m0_re_rom[23] = 128;
    assign twf_m0_im_rom[23] = 0;
    assign twf_m0_re_rom[24] = 128;
    assign twf_m0_im_rom[24] = 0;
    assign twf_m0_re_rom[25] = 128;
    assign twf_m0_im_rom[25] = 0;
    assign twf_m0_re_rom[26] = 128;
    assign twf_m0_im_rom[26] = 0;
    assign twf_m0_re_rom[27] = 128;
    assign twf_m0_im_rom[27] = 0;
    assign twf_m0_re_rom[28] = 128;
    assign twf_m0_im_rom[28] = 0;
    assign twf_m0_re_rom[29] = 128;
    assign twf_m0_im_rom[29] = 0;
    assign twf_m0_re_rom[30] = 128;
    assign twf_m0_im_rom[30] = 0;
    assign twf_m0_re_rom[31] = 128;
    assign twf_m0_im_rom[31] = 0;
    assign twf_m0_re_rom[32] = 128;
    assign twf_m0_im_rom[32] = 0;
    assign twf_m0_re_rom[33] = 128;
    assign twf_m0_im_rom[33] = 0;
    assign twf_m0_re_rom[34] = 128;
    assign twf_m0_im_rom[34] = 0;
    assign twf_m0_re_rom[35] = 128;
    assign twf_m0_im_rom[35] = 0;
    assign twf_m0_re_rom[36] = 128;
    assign twf_m0_im_rom[36] = 0;
    assign twf_m0_re_rom[37] = 128;
    assign twf_m0_im_rom[37] = 0;
    assign twf_m0_re_rom[38] = 128;
    assign twf_m0_im_rom[38] = 0;
    assign twf_m0_re_rom[39] = 128;
    assign twf_m0_im_rom[39] = 0;
    assign twf_m0_re_rom[40] = 128;
    assign twf_m0_im_rom[40] = 0;
    assign twf_m0_re_rom[41] = 128;
    assign twf_m0_im_rom[41] = 0;
    assign twf_m0_re_rom[42] = 128;
    assign twf_m0_im_rom[42] = 0;
    assign twf_m0_re_rom[43] = 128;
    assign twf_m0_im_rom[43] = 0;
    assign twf_m0_re_rom[44] = 128;
    assign twf_m0_im_rom[44] = 0;
    assign twf_m0_re_rom[45] = 128;
    assign twf_m0_im_rom[45] = 0;
    assign twf_m0_re_rom[46] = 128;
    assign twf_m0_im_rom[46] = 0;
    assign twf_m0_re_rom[47] = 128;
    assign twf_m0_im_rom[47] = 0;
    assign twf_m0_re_rom[48] = 128;
    assign twf_m0_im_rom[48] = 0;
    assign twf_m0_re_rom[49] = 128;
    assign twf_m0_im_rom[49] = 0;
    assign twf_m0_re_rom[50] = 128;
    assign twf_m0_im_rom[50] = 0;
    assign twf_m0_re_rom[51] = 128;
    assign twf_m0_im_rom[51] = 0;
    assign twf_m0_re_rom[52] = 128;
    assign twf_m0_im_rom[52] = 0;
    assign twf_m0_re_rom[53] = 128;
    assign twf_m0_im_rom[53] = 0;
    assign twf_m0_re_rom[54] = 128;
    assign twf_m0_im_rom[54] = 0;
    assign twf_m0_re_rom[55] = 128;
    assign twf_m0_im_rom[55] = 0;
    assign twf_m0_re_rom[56] = 128;
    assign twf_m0_im_rom[56] = 0;
    assign twf_m0_re_rom[57] = 128;
    assign twf_m0_im_rom[57] = 0;
    assign twf_m0_re_rom[58] = 128;
    assign twf_m0_im_rom[58] = 0;
    assign twf_m0_re_rom[59] = 128;
    assign twf_m0_im_rom[59] = 0;
    assign twf_m0_re_rom[60] = 128;
    assign twf_m0_im_rom[60] = 0;
    assign twf_m0_re_rom[61] = 128;
    assign twf_m0_im_rom[61] = 0;
    assign twf_m0_re_rom[62] = 128;
    assign twf_m0_im_rom[62] = 0;
    assign twf_m0_re_rom[63] = 128;
    assign twf_m0_im_rom[63] = 0;
    assign twf_m0_re_rom[64] = 128;
    assign twf_m0_im_rom[64] = 0;
    assign twf_m0_re_rom[65] = 128;
    assign twf_m0_im_rom[65] = -6;
    assign twf_m0_re_rom[66] = 127;
    assign twf_m0_im_rom[66] = -13;
    assign twf_m0_re_rom[67] = 127;
    assign twf_m0_im_rom[67] = -19;
    assign twf_m0_re_rom[68] = 126;
    assign twf_m0_im_rom[68] = -25;
    assign twf_m0_re_rom[69] = 124;
    assign twf_m0_im_rom[69] = -31;
    assign twf_m0_re_rom[70] = 122;
    assign twf_m0_im_rom[70] = -37;
    assign twf_m0_re_rom[71] = 121;
    assign twf_m0_im_rom[71] = -43;
    assign twf_m0_re_rom[72] = 118;
    assign twf_m0_im_rom[72] = -49;
    assign twf_m0_re_rom[73] = 116;
    assign twf_m0_im_rom[73] = -55;
    assign twf_m0_re_rom[74] = 113;
    assign twf_m0_im_rom[74] = -60;
    assign twf_m0_re_rom[75] = 110;
    assign twf_m0_im_rom[75] = -66;
    assign twf_m0_re_rom[76] = 106;
    assign twf_m0_im_rom[76] = -71;
    assign twf_m0_re_rom[77] = 103;
    assign twf_m0_im_rom[77] = -76;
    assign twf_m0_re_rom[78] = 99;
    assign twf_m0_im_rom[78] = -81;
    assign twf_m0_re_rom[79] = 95;
    assign twf_m0_im_rom[79] = -86;
    assign twf_m0_re_rom[80] = 91;
    assign twf_m0_im_rom[80] = -91;
    assign twf_m0_re_rom[81] = 86;
    assign twf_m0_im_rom[81] = -95;
    assign twf_m0_re_rom[82] = 81;
    assign twf_m0_im_rom[82] = -99;
    assign twf_m0_re_rom[83] = 76;
    assign twf_m0_im_rom[83] = -103;
    assign twf_m0_re_rom[84] = 71;
    assign twf_m0_im_rom[84] = -106;
    assign twf_m0_re_rom[85] = 66;
    assign twf_m0_im_rom[85] = -110;
    assign twf_m0_re_rom[86] = 60;
    assign twf_m0_im_rom[86] = -113;
    assign twf_m0_re_rom[87] = 55;
    assign twf_m0_im_rom[87] = -116;
    assign twf_m0_re_rom[88] = 49;
    assign twf_m0_im_rom[88] = -118;
    assign twf_m0_re_rom[89] = 43;
    assign twf_m0_im_rom[89] = -121;
    assign twf_m0_re_rom[90] = 37;
    assign twf_m0_im_rom[90] = -122;
    assign twf_m0_re_rom[91] = 31;
    assign twf_m0_im_rom[91] = -124;
    assign twf_m0_re_rom[92] = 25;
    assign twf_m0_im_rom[92] = -126;
    assign twf_m0_re_rom[93] = 19;
    assign twf_m0_im_rom[93] = -127;
    assign twf_m0_re_rom[94] = 13;
    assign twf_m0_im_rom[94] = -127;
    assign twf_m0_re_rom[95] = 6;
    assign twf_m0_im_rom[95] = -128;
    assign twf_m0_re_rom[96] = 0;
    assign twf_m0_im_rom[96] = -128;
    assign twf_m0_re_rom[97] = -6;
    assign twf_m0_im_rom[97] = -128;
    assign twf_m0_re_rom[98] = -13;
    assign twf_m0_im_rom[98] = -127;
    assign twf_m0_re_rom[99] = -19;
    assign twf_m0_im_rom[99] = -127;
    assign twf_m0_re_rom[100] = -25;
    assign twf_m0_im_rom[100] = -126;
    assign twf_m0_re_rom[101] = -31;
    assign twf_m0_im_rom[101] = -124;
    assign twf_m0_re_rom[102] = -37;
    assign twf_m0_im_rom[102] = -122;
    assign twf_m0_re_rom[103] = -43;
    assign twf_m0_im_rom[103] = -121;
    assign twf_m0_re_rom[104] = -49;
    assign twf_m0_im_rom[104] = -118;
    assign twf_m0_re_rom[105] = -55;
    assign twf_m0_im_rom[105] = -116;
    assign twf_m0_re_rom[106] = -60;
    assign twf_m0_im_rom[106] = -113;
    assign twf_m0_re_rom[107] = -66;
    assign twf_m0_im_rom[107] = -110;
    assign twf_m0_re_rom[108] = -71;
    assign twf_m0_im_rom[108] = -106;
    assign twf_m0_re_rom[109] = -76;
    assign twf_m0_im_rom[109] = -103;
    assign twf_m0_re_rom[110] = -81;
    assign twf_m0_im_rom[110] = -99;
    assign twf_m0_re_rom[111] = -86;
    assign twf_m0_im_rom[111] = -95;
    assign twf_m0_re_rom[112] = -91;
    assign twf_m0_im_rom[112] = -91;
    assign twf_m0_re_rom[113] = -95;
    assign twf_m0_im_rom[113] = -86;
    assign twf_m0_re_rom[114] = -99;
    assign twf_m0_im_rom[114] = -81;
    assign twf_m0_re_rom[115] = -103;
    assign twf_m0_im_rom[115] = -76;
    assign twf_m0_re_rom[116] = -106;
    assign twf_m0_im_rom[116] = -71;
    assign twf_m0_re_rom[117] = -110;
    assign twf_m0_im_rom[117] = -66;
    assign twf_m0_re_rom[118] = -113;
    assign twf_m0_im_rom[118] = -60;
    assign twf_m0_re_rom[119] = -116;
    assign twf_m0_im_rom[119] = -55;
    assign twf_m0_re_rom[120] = -118;
    assign twf_m0_im_rom[120] = -49;
    assign twf_m0_re_rom[121] = -121;
    assign twf_m0_im_rom[121] = -43;
    assign twf_m0_re_rom[122] = -122;
    assign twf_m0_im_rom[122] = -37;
    assign twf_m0_re_rom[123] = -124;
    assign twf_m0_im_rom[123] = -31;
    assign twf_m0_re_rom[124] = -126;
    assign twf_m0_im_rom[124] = -25;
    assign twf_m0_re_rom[125] = -127;
    assign twf_m0_im_rom[125] = -19;
    assign twf_m0_re_rom[126] = -127;
    assign twf_m0_im_rom[126] = -13;
    assign twf_m0_re_rom[127] = -128;
    assign twf_m0_im_rom[127] = -6;
    assign twf_m0_re_rom[128] = 128;
    assign twf_m0_im_rom[128] = 0;
    assign twf_m0_re_rom[129] = 128;
    assign twf_m0_im_rom[129] = -3;
    assign twf_m0_re_rom[130] = 128;
    assign twf_m0_im_rom[130] = -6;
    assign twf_m0_re_rom[131] = 128;
    assign twf_m0_im_rom[131] = -9;
    assign twf_m0_re_rom[132] = 127;
    assign twf_m0_im_rom[132] = -13;
    assign twf_m0_re_rom[133] = 127;
    assign twf_m0_im_rom[133] = -16;
    assign twf_m0_re_rom[134] = 127;
    assign twf_m0_im_rom[134] = -19;
    assign twf_m0_re_rom[135] = 126;
    assign twf_m0_im_rom[135] = -22;
    assign twf_m0_re_rom[136] = 126;
    assign twf_m0_im_rom[136] = -25;
    assign twf_m0_re_rom[137] = 125;
    assign twf_m0_im_rom[137] = -28;
    assign twf_m0_re_rom[138] = 124;
    assign twf_m0_im_rom[138] = -31;
    assign twf_m0_re_rom[139] = 123;
    assign twf_m0_im_rom[139] = -34;
    assign twf_m0_re_rom[140] = 122;
    assign twf_m0_im_rom[140] = -37;
    assign twf_m0_re_rom[141] = 122;
    assign twf_m0_im_rom[141] = -40;
    assign twf_m0_re_rom[142] = 121;
    assign twf_m0_im_rom[142] = -43;
    assign twf_m0_re_rom[143] = 119;
    assign twf_m0_im_rom[143] = -46;
    assign twf_m0_re_rom[144] = 118;
    assign twf_m0_im_rom[144] = -49;
    assign twf_m0_re_rom[145] = 117;
    assign twf_m0_im_rom[145] = -52;
    assign twf_m0_re_rom[146] = 116;
    assign twf_m0_im_rom[146] = -55;
    assign twf_m0_re_rom[147] = 114;
    assign twf_m0_im_rom[147] = -58;
    assign twf_m0_re_rom[148] = 113;
    assign twf_m0_im_rom[148] = -60;
    assign twf_m0_re_rom[149] = 111;
    assign twf_m0_im_rom[149] = -63;
    assign twf_m0_re_rom[150] = 110;
    assign twf_m0_im_rom[150] = -66;
    assign twf_m0_re_rom[151] = 108;
    assign twf_m0_im_rom[151] = -68;
    assign twf_m0_re_rom[152] = 106;
    assign twf_m0_im_rom[152] = -71;
    assign twf_m0_re_rom[153] = 105;
    assign twf_m0_im_rom[153] = -74;
    assign twf_m0_re_rom[154] = 103;
    assign twf_m0_im_rom[154] = -76;
    assign twf_m0_re_rom[155] = 101;
    assign twf_m0_im_rom[155] = -79;
    assign twf_m0_re_rom[156] = 99;
    assign twf_m0_im_rom[156] = -81;
    assign twf_m0_re_rom[157] = 97;
    assign twf_m0_im_rom[157] = -84;
    assign twf_m0_re_rom[158] = 95;
    assign twf_m0_im_rom[158] = -86;
    assign twf_m0_re_rom[159] = 93;
    assign twf_m0_im_rom[159] = -88;
    assign twf_m0_re_rom[160] = 91;
    assign twf_m0_im_rom[160] = -91;
    assign twf_m0_re_rom[161] = 88;
    assign twf_m0_im_rom[161] = -93;
    assign twf_m0_re_rom[162] = 86;
    assign twf_m0_im_rom[162] = -95;
    assign twf_m0_re_rom[163] = 84;
    assign twf_m0_im_rom[163] = -97;
    assign twf_m0_re_rom[164] = 81;
    assign twf_m0_im_rom[164] = -99;
    assign twf_m0_re_rom[165] = 79;
    assign twf_m0_im_rom[165] = -101;
    assign twf_m0_re_rom[166] = 76;
    assign twf_m0_im_rom[166] = -103;
    assign twf_m0_re_rom[167] = 74;
    assign twf_m0_im_rom[167] = -105;
    assign twf_m0_re_rom[168] = 71;
    assign twf_m0_im_rom[168] = -106;
    assign twf_m0_re_rom[169] = 68;
    assign twf_m0_im_rom[169] = -108;
    assign twf_m0_re_rom[170] = 66;
    assign twf_m0_im_rom[170] = -110;
    assign twf_m0_re_rom[171] = 63;
    assign twf_m0_im_rom[171] = -111;
    assign twf_m0_re_rom[172] = 60;
    assign twf_m0_im_rom[172] = -113;
    assign twf_m0_re_rom[173] = 58;
    assign twf_m0_im_rom[173] = -114;
    assign twf_m0_re_rom[174] = 55;
    assign twf_m0_im_rom[174] = -116;
    assign twf_m0_re_rom[175] = 52;
    assign twf_m0_im_rom[175] = -117;
    assign twf_m0_re_rom[176] = 49;
    assign twf_m0_im_rom[176] = -118;
    assign twf_m0_re_rom[177] = 46;
    assign twf_m0_im_rom[177] = -119;
    assign twf_m0_re_rom[178] = 43;
    assign twf_m0_im_rom[178] = -121;
    assign twf_m0_re_rom[179] = 40;
    assign twf_m0_im_rom[179] = -122;
    assign twf_m0_re_rom[180] = 37;
    assign twf_m0_im_rom[180] = -122;
    assign twf_m0_re_rom[181] = 34;
    assign twf_m0_im_rom[181] = -123;
    assign twf_m0_re_rom[182] = 31;
    assign twf_m0_im_rom[182] = -124;
    assign twf_m0_re_rom[183] = 28;
    assign twf_m0_im_rom[183] = -125;
    assign twf_m0_re_rom[184] = 25;
    assign twf_m0_im_rom[184] = -126;
    assign twf_m0_re_rom[185] = 22;
    assign twf_m0_im_rom[185] = -126;
    assign twf_m0_re_rom[186] = 19;
    assign twf_m0_im_rom[186] = -127;
    assign twf_m0_re_rom[187] = 16;
    assign twf_m0_im_rom[187] = -127;
    assign twf_m0_re_rom[188] = 13;
    assign twf_m0_im_rom[188] = -127;
    assign twf_m0_re_rom[189] = 9;
    assign twf_m0_im_rom[189] = -128;
    assign twf_m0_re_rom[190] = 6;
    assign twf_m0_im_rom[190] = -128;
    assign twf_m0_re_rom[191] = 3;
    assign twf_m0_im_rom[191] = -128;
    assign twf_m0_re_rom[192] = 128;
    assign twf_m0_im_rom[192] = 0;
    assign twf_m0_re_rom[193] = 128;
    assign twf_m0_im_rom[193] = -9;
    assign twf_m0_re_rom[194] = 127;
    assign twf_m0_im_rom[194] = -19;
    assign twf_m0_re_rom[195] = 125;
    assign twf_m0_im_rom[195] = -28;
    assign twf_m0_re_rom[196] = 122;
    assign twf_m0_im_rom[196] = -37;
    assign twf_m0_re_rom[197] = 119;
    assign twf_m0_im_rom[197] = -46;
    assign twf_m0_re_rom[198] = 116;
    assign twf_m0_im_rom[198] = -55;
    assign twf_m0_re_rom[199] = 111;
    assign twf_m0_im_rom[199] = -63;
    assign twf_m0_re_rom[200] = 106;
    assign twf_m0_im_rom[200] = -71;
    assign twf_m0_re_rom[201] = 101;
    assign twf_m0_im_rom[201] = -79;
    assign twf_m0_re_rom[202] = 95;
    assign twf_m0_im_rom[202] = -86;
    assign twf_m0_re_rom[203] = 88;
    assign twf_m0_im_rom[203] = -93;
    assign twf_m0_re_rom[204] = 81;
    assign twf_m0_im_rom[204] = -99;
    assign twf_m0_re_rom[205] = 74;
    assign twf_m0_im_rom[205] = -105;
    assign twf_m0_re_rom[206] = 66;
    assign twf_m0_im_rom[206] = -110;
    assign twf_m0_re_rom[207] = 58;
    assign twf_m0_im_rom[207] = -114;
    assign twf_m0_re_rom[208] = 49;
    assign twf_m0_im_rom[208] = -118;
    assign twf_m0_re_rom[209] = 40;
    assign twf_m0_im_rom[209] = -122;
    assign twf_m0_re_rom[210] = 31;
    assign twf_m0_im_rom[210] = -124;
    assign twf_m0_re_rom[211] = 22;
    assign twf_m0_im_rom[211] = -126;
    assign twf_m0_re_rom[212] = 13;
    assign twf_m0_im_rom[212] = -127;
    assign twf_m0_re_rom[213] = 3;
    assign twf_m0_im_rom[213] = -128;
    assign twf_m0_re_rom[214] = -6;
    assign twf_m0_im_rom[214] = -128;
    assign twf_m0_re_rom[215] = -16;
    assign twf_m0_im_rom[215] = -127;
    assign twf_m0_re_rom[216] = -25;
    assign twf_m0_im_rom[216] = -126;
    assign twf_m0_re_rom[217] = -34;
    assign twf_m0_im_rom[217] = -123;
    assign twf_m0_re_rom[218] = -43;
    assign twf_m0_im_rom[218] = -121;
    assign twf_m0_re_rom[219] = -52;
    assign twf_m0_im_rom[219] = -117;
    assign twf_m0_re_rom[220] = -60;
    assign twf_m0_im_rom[220] = -113;
    assign twf_m0_re_rom[221] = -68;
    assign twf_m0_im_rom[221] = -108;
    assign twf_m0_re_rom[222] = -76;
    assign twf_m0_im_rom[222] = -103;
    assign twf_m0_re_rom[223] = -84;
    assign twf_m0_im_rom[223] = -97;
    assign twf_m0_re_rom[224] = -91;
    assign twf_m0_im_rom[224] = -91;
    assign twf_m0_re_rom[225] = -97;
    assign twf_m0_im_rom[225] = -84;
    assign twf_m0_re_rom[226] = -103;
    assign twf_m0_im_rom[226] = -76;
    assign twf_m0_re_rom[227] = -108;
    assign twf_m0_im_rom[227] = -68;
    assign twf_m0_re_rom[228] = -113;
    assign twf_m0_im_rom[228] = -60;
    assign twf_m0_re_rom[229] = -117;
    assign twf_m0_im_rom[229] = -52;
    assign twf_m0_re_rom[230] = -121;
    assign twf_m0_im_rom[230] = -43;
    assign twf_m0_re_rom[231] = -123;
    assign twf_m0_im_rom[231] = -34;
    assign twf_m0_re_rom[232] = -126;
    assign twf_m0_im_rom[232] = -25;
    assign twf_m0_re_rom[233] = -127;
    assign twf_m0_im_rom[233] = -16;
    assign twf_m0_re_rom[234] = -128;
    assign twf_m0_im_rom[234] = -6;
    assign twf_m0_re_rom[235] = -128;
    assign twf_m0_im_rom[235] = 3;
    assign twf_m0_re_rom[236] = -127;
    assign twf_m0_im_rom[236] = 13;
    assign twf_m0_re_rom[237] = -126;
    assign twf_m0_im_rom[237] = 22;
    assign twf_m0_re_rom[238] = -124;
    assign twf_m0_im_rom[238] = 31;
    assign twf_m0_re_rom[239] = -122;
    assign twf_m0_im_rom[239] = 40;
    assign twf_m0_re_rom[240] = -118;
    assign twf_m0_im_rom[240] = 49;
    assign twf_m0_re_rom[241] = -114;
    assign twf_m0_im_rom[241] = 58;
    assign twf_m0_re_rom[242] = -110;
    assign twf_m0_im_rom[242] = 66;
    assign twf_m0_re_rom[243] = -105;
    assign twf_m0_im_rom[243] = 74;
    assign twf_m0_re_rom[244] = -99;
    assign twf_m0_im_rom[244] = 81;
    assign twf_m0_re_rom[245] = -93;
    assign twf_m0_im_rom[245] = 88;
    assign twf_m0_re_rom[246] = -86;
    assign twf_m0_im_rom[246] = 95;
    assign twf_m0_re_rom[247] = -79;
    assign twf_m0_im_rom[247] = 101;
    assign twf_m0_re_rom[248] = -71;
    assign twf_m0_im_rom[248] = 106;
    assign twf_m0_re_rom[249] = -63;
    assign twf_m0_im_rom[249] = 111;
    assign twf_m0_re_rom[250] = -55;
    assign twf_m0_im_rom[250] = 116;
    assign twf_m0_re_rom[251] = -46;
    assign twf_m0_im_rom[251] = 119;
    assign twf_m0_re_rom[252] = -37;
    assign twf_m0_im_rom[252] = 122;
    assign twf_m0_re_rom[253] = -28;
    assign twf_m0_im_rom[253] = 125;
    assign twf_m0_re_rom[254] = -19;
    assign twf_m0_im_rom[254] = 127;
    assign twf_m0_re_rom[255] = -9;
    assign twf_m0_im_rom[255] = 128;
    assign twf_m0_re_rom[256] = 128;
    assign twf_m0_im_rom[256] = 0;
    assign twf_m0_re_rom[257] = 128;
    assign twf_m0_im_rom[257] = -2;
    assign twf_m0_re_rom[258] = 128;
    assign twf_m0_im_rom[258] = -3;
    assign twf_m0_re_rom[259] = 128;
    assign twf_m0_im_rom[259] = -5;
    assign twf_m0_re_rom[260] = 128;
    assign twf_m0_im_rom[260] = -6;
    assign twf_m0_re_rom[261] = 128;
    assign twf_m0_im_rom[261] = -8;
    assign twf_m0_re_rom[262] = 128;
    assign twf_m0_im_rom[262] = -9;
    assign twf_m0_re_rom[263] = 128;
    assign twf_m0_im_rom[263] = -11;
    assign twf_m0_re_rom[264] = 127;
    assign twf_m0_im_rom[264] = -13;
    assign twf_m0_re_rom[265] = 127;
    assign twf_m0_im_rom[265] = -14;
    assign twf_m0_re_rom[266] = 127;
    assign twf_m0_im_rom[266] = -16;
    assign twf_m0_re_rom[267] = 127;
    assign twf_m0_im_rom[267] = -17;
    assign twf_m0_re_rom[268] = 127;
    assign twf_m0_im_rom[268] = -19;
    assign twf_m0_re_rom[269] = 126;
    assign twf_m0_im_rom[269] = -20;
    assign twf_m0_re_rom[270] = 126;
    assign twf_m0_im_rom[270] = -22;
    assign twf_m0_re_rom[271] = 126;
    assign twf_m0_im_rom[271] = -23;
    assign twf_m0_re_rom[272] = 126;
    assign twf_m0_im_rom[272] = -25;
    assign twf_m0_re_rom[273] = 125;
    assign twf_m0_im_rom[273] = -27;
    assign twf_m0_re_rom[274] = 125;
    assign twf_m0_im_rom[274] = -28;
    assign twf_m0_re_rom[275] = 125;
    assign twf_m0_im_rom[275] = -30;
    assign twf_m0_re_rom[276] = 124;
    assign twf_m0_im_rom[276] = -31;
    assign twf_m0_re_rom[277] = 124;
    assign twf_m0_im_rom[277] = -33;
    assign twf_m0_re_rom[278] = 123;
    assign twf_m0_im_rom[278] = -34;
    assign twf_m0_re_rom[279] = 123;
    assign twf_m0_im_rom[279] = -36;
    assign twf_m0_re_rom[280] = 122;
    assign twf_m0_im_rom[280] = -37;
    assign twf_m0_re_rom[281] = 122;
    assign twf_m0_im_rom[281] = -39;
    assign twf_m0_re_rom[282] = 122;
    assign twf_m0_im_rom[282] = -40;
    assign twf_m0_re_rom[283] = 121;
    assign twf_m0_im_rom[283] = -42;
    assign twf_m0_re_rom[284] = 121;
    assign twf_m0_im_rom[284] = -43;
    assign twf_m0_re_rom[285] = 120;
    assign twf_m0_im_rom[285] = -45;
    assign twf_m0_re_rom[286] = 119;
    assign twf_m0_im_rom[286] = -46;
    assign twf_m0_re_rom[287] = 119;
    assign twf_m0_im_rom[287] = -48;
    assign twf_m0_re_rom[288] = 118;
    assign twf_m0_im_rom[288] = -49;
    assign twf_m0_re_rom[289] = 118;
    assign twf_m0_im_rom[289] = -50;
    assign twf_m0_re_rom[290] = 117;
    assign twf_m0_im_rom[290] = -52;
    assign twf_m0_re_rom[291] = 116;
    assign twf_m0_im_rom[291] = -53;
    assign twf_m0_re_rom[292] = 116;
    assign twf_m0_im_rom[292] = -55;
    assign twf_m0_re_rom[293] = 115;
    assign twf_m0_im_rom[293] = -56;
    assign twf_m0_re_rom[294] = 114;
    assign twf_m0_im_rom[294] = -58;
    assign twf_m0_re_rom[295] = 114;
    assign twf_m0_im_rom[295] = -59;
    assign twf_m0_re_rom[296] = 113;
    assign twf_m0_im_rom[296] = -60;
    assign twf_m0_re_rom[297] = 112;
    assign twf_m0_im_rom[297] = -62;
    assign twf_m0_re_rom[298] = 111;
    assign twf_m0_im_rom[298] = -63;
    assign twf_m0_re_rom[299] = 111;
    assign twf_m0_im_rom[299] = -64;
    assign twf_m0_re_rom[300] = 110;
    assign twf_m0_im_rom[300] = -66;
    assign twf_m0_re_rom[301] = 109;
    assign twf_m0_im_rom[301] = -67;
    assign twf_m0_re_rom[302] = 108;
    assign twf_m0_im_rom[302] = -68;
    assign twf_m0_re_rom[303] = 107;
    assign twf_m0_im_rom[303] = -70;
    assign twf_m0_re_rom[304] = 106;
    assign twf_m0_im_rom[304] = -71;
    assign twf_m0_re_rom[305] = 106;
    assign twf_m0_im_rom[305] = -72;
    assign twf_m0_re_rom[306] = 105;
    assign twf_m0_im_rom[306] = -74;
    assign twf_m0_re_rom[307] = 104;
    assign twf_m0_im_rom[307] = -75;
    assign twf_m0_re_rom[308] = 103;
    assign twf_m0_im_rom[308] = -76;
    assign twf_m0_re_rom[309] = 102;
    assign twf_m0_im_rom[309] = -78;
    assign twf_m0_re_rom[310] = 101;
    assign twf_m0_im_rom[310] = -79;
    assign twf_m0_re_rom[311] = 100;
    assign twf_m0_im_rom[311] = -80;
    assign twf_m0_re_rom[312] = 99;
    assign twf_m0_im_rom[312] = -81;
    assign twf_m0_re_rom[313] = 98;
    assign twf_m0_im_rom[313] = -82;
    assign twf_m0_re_rom[314] = 97;
    assign twf_m0_im_rom[314] = -84;
    assign twf_m0_re_rom[315] = 96;
    assign twf_m0_im_rom[315] = -85;
    assign twf_m0_re_rom[316] = 95;
    assign twf_m0_im_rom[316] = -86;
    assign twf_m0_re_rom[317] = 94;
    assign twf_m0_im_rom[317] = -87;
    assign twf_m0_re_rom[318] = 93;
    assign twf_m0_im_rom[318] = -88;
    assign twf_m0_re_rom[319] = 92;
    assign twf_m0_im_rom[319] = -89;
    assign twf_m0_re_rom[320] = 128;
    assign twf_m0_im_rom[320] = 0;
    assign twf_m0_re_rom[321] = 128;
    assign twf_m0_im_rom[321] = -8;
    assign twf_m0_re_rom[322] = 127;
    assign twf_m0_im_rom[322] = -16;
    assign twf_m0_re_rom[323] = 126;
    assign twf_m0_im_rom[323] = -23;
    assign twf_m0_re_rom[324] = 124;
    assign twf_m0_im_rom[324] = -31;
    assign twf_m0_re_rom[325] = 122;
    assign twf_m0_im_rom[325] = -39;
    assign twf_m0_re_rom[326] = 119;
    assign twf_m0_im_rom[326] = -46;
    assign twf_m0_re_rom[327] = 116;
    assign twf_m0_im_rom[327] = -53;
    assign twf_m0_re_rom[328] = 113;
    assign twf_m0_im_rom[328] = -60;
    assign twf_m0_re_rom[329] = 109;
    assign twf_m0_im_rom[329] = -67;
    assign twf_m0_re_rom[330] = 105;
    assign twf_m0_im_rom[330] = -74;
    assign twf_m0_re_rom[331] = 100;
    assign twf_m0_im_rom[331] = -80;
    assign twf_m0_re_rom[332] = 95;
    assign twf_m0_im_rom[332] = -86;
    assign twf_m0_re_rom[333] = 89;
    assign twf_m0_im_rom[333] = -92;
    assign twf_m0_re_rom[334] = 84;
    assign twf_m0_im_rom[334] = -97;
    assign twf_m0_re_rom[335] = 78;
    assign twf_m0_im_rom[335] = -102;
    assign twf_m0_re_rom[336] = 71;
    assign twf_m0_im_rom[336] = -106;
    assign twf_m0_re_rom[337] = 64;
    assign twf_m0_im_rom[337] = -111;
    assign twf_m0_re_rom[338] = 58;
    assign twf_m0_im_rom[338] = -114;
    assign twf_m0_re_rom[339] = 50;
    assign twf_m0_im_rom[339] = -118;
    assign twf_m0_re_rom[340] = 43;
    assign twf_m0_im_rom[340] = -121;
    assign twf_m0_re_rom[341] = 36;
    assign twf_m0_im_rom[341] = -123;
    assign twf_m0_re_rom[342] = 28;
    assign twf_m0_im_rom[342] = -125;
    assign twf_m0_re_rom[343] = 20;
    assign twf_m0_im_rom[343] = -126;
    assign twf_m0_re_rom[344] = 13;
    assign twf_m0_im_rom[344] = -127;
    assign twf_m0_re_rom[345] = 5;
    assign twf_m0_im_rom[345] = -128;
    assign twf_m0_re_rom[346] = -3;
    assign twf_m0_im_rom[346] = -128;
    assign twf_m0_re_rom[347] = -11;
    assign twf_m0_im_rom[347] = -128;
    assign twf_m0_re_rom[348] = -19;
    assign twf_m0_im_rom[348] = -127;
    assign twf_m0_re_rom[349] = -27;
    assign twf_m0_im_rom[349] = -125;
    assign twf_m0_re_rom[350] = -34;
    assign twf_m0_im_rom[350] = -123;
    assign twf_m0_re_rom[351] = -42;
    assign twf_m0_im_rom[351] = -121;
    assign twf_m0_re_rom[352] = -49;
    assign twf_m0_im_rom[352] = -118;
    assign twf_m0_re_rom[353] = -56;
    assign twf_m0_im_rom[353] = -115;
    assign twf_m0_re_rom[354] = -63;
    assign twf_m0_im_rom[354] = -111;
    assign twf_m0_re_rom[355] = -70;
    assign twf_m0_im_rom[355] = -107;
    assign twf_m0_re_rom[356] = -76;
    assign twf_m0_im_rom[356] = -103;
    assign twf_m0_re_rom[357] = -82;
    assign twf_m0_im_rom[357] = -98;
    assign twf_m0_re_rom[358] = -88;
    assign twf_m0_im_rom[358] = -93;
    assign twf_m0_re_rom[359] = -94;
    assign twf_m0_im_rom[359] = -87;
    assign twf_m0_re_rom[360] = -99;
    assign twf_m0_im_rom[360] = -81;
    assign twf_m0_re_rom[361] = -104;
    assign twf_m0_im_rom[361] = -75;
    assign twf_m0_re_rom[362] = -108;
    assign twf_m0_im_rom[362] = -68;
    assign twf_m0_re_rom[363] = -112;
    assign twf_m0_im_rom[363] = -62;
    assign twf_m0_re_rom[364] = -116;
    assign twf_m0_im_rom[364] = -55;
    assign twf_m0_re_rom[365] = -119;
    assign twf_m0_im_rom[365] = -48;
    assign twf_m0_re_rom[366] = -122;
    assign twf_m0_im_rom[366] = -40;
    assign twf_m0_re_rom[367] = -124;
    assign twf_m0_im_rom[367] = -33;
    assign twf_m0_re_rom[368] = -126;
    assign twf_m0_im_rom[368] = -25;
    assign twf_m0_re_rom[369] = -127;
    assign twf_m0_im_rom[369] = -17;
    assign twf_m0_re_rom[370] = -128;
    assign twf_m0_im_rom[370] = -9;
    assign twf_m0_re_rom[371] = -128;
    assign twf_m0_im_rom[371] = -2;
    assign twf_m0_re_rom[372] = -128;
    assign twf_m0_im_rom[372] = 6;
    assign twf_m0_re_rom[373] = -127;
    assign twf_m0_im_rom[373] = 14;
    assign twf_m0_re_rom[374] = -126;
    assign twf_m0_im_rom[374] = 22;
    assign twf_m0_re_rom[375] = -125;
    assign twf_m0_im_rom[375] = 30;
    assign twf_m0_re_rom[376] = -122;
    assign twf_m0_im_rom[376] = 37;
    assign twf_m0_re_rom[377] = -120;
    assign twf_m0_im_rom[377] = 45;
    assign twf_m0_re_rom[378] = -117;
    assign twf_m0_im_rom[378] = 52;
    assign twf_m0_re_rom[379] = -114;
    assign twf_m0_im_rom[379] = 59;
    assign twf_m0_re_rom[380] = -110;
    assign twf_m0_im_rom[380] = 66;
    assign twf_m0_re_rom[381] = -106;
    assign twf_m0_im_rom[381] = 72;
    assign twf_m0_re_rom[382] = -101;
    assign twf_m0_im_rom[382] = 79;
    assign twf_m0_re_rom[383] = -96;
    assign twf_m0_im_rom[383] = 85;
    assign twf_m0_re_rom[384] = 128;
    assign twf_m0_im_rom[384] = 0;
    assign twf_m0_re_rom[385] = 128;
    assign twf_m0_im_rom[385] = -5;
    assign twf_m0_re_rom[386] = 128;
    assign twf_m0_im_rom[386] = -9;
    assign twf_m0_re_rom[387] = 127;
    assign twf_m0_im_rom[387] = -14;
    assign twf_m0_re_rom[388] = 127;
    assign twf_m0_im_rom[388] = -19;
    assign twf_m0_re_rom[389] = 126;
    assign twf_m0_im_rom[389] = -23;
    assign twf_m0_re_rom[390] = 125;
    assign twf_m0_im_rom[390] = -28;
    assign twf_m0_re_rom[391] = 124;
    assign twf_m0_im_rom[391] = -33;
    assign twf_m0_re_rom[392] = 122;
    assign twf_m0_im_rom[392] = -37;
    assign twf_m0_re_rom[393] = 121;
    assign twf_m0_im_rom[393] = -42;
    assign twf_m0_re_rom[394] = 119;
    assign twf_m0_im_rom[394] = -46;
    assign twf_m0_re_rom[395] = 118;
    assign twf_m0_im_rom[395] = -50;
    assign twf_m0_re_rom[396] = 116;
    assign twf_m0_im_rom[396] = -55;
    assign twf_m0_re_rom[397] = 114;
    assign twf_m0_im_rom[397] = -59;
    assign twf_m0_re_rom[398] = 111;
    assign twf_m0_im_rom[398] = -63;
    assign twf_m0_re_rom[399] = 109;
    assign twf_m0_im_rom[399] = -67;
    assign twf_m0_re_rom[400] = 106;
    assign twf_m0_im_rom[400] = -71;
    assign twf_m0_re_rom[401] = 104;
    assign twf_m0_im_rom[401] = -75;
    assign twf_m0_re_rom[402] = 101;
    assign twf_m0_im_rom[402] = -79;
    assign twf_m0_re_rom[403] = 98;
    assign twf_m0_im_rom[403] = -82;
    assign twf_m0_re_rom[404] = 95;
    assign twf_m0_im_rom[404] = -86;
    assign twf_m0_re_rom[405] = 92;
    assign twf_m0_im_rom[405] = -89;
    assign twf_m0_re_rom[406] = 88;
    assign twf_m0_im_rom[406] = -93;
    assign twf_m0_re_rom[407] = 85;
    assign twf_m0_im_rom[407] = -96;
    assign twf_m0_re_rom[408] = 81;
    assign twf_m0_im_rom[408] = -99;
    assign twf_m0_re_rom[409] = 78;
    assign twf_m0_im_rom[409] = -102;
    assign twf_m0_re_rom[410] = 74;
    assign twf_m0_im_rom[410] = -105;
    assign twf_m0_re_rom[411] = 70;
    assign twf_m0_im_rom[411] = -107;
    assign twf_m0_re_rom[412] = 66;
    assign twf_m0_im_rom[412] = -110;
    assign twf_m0_re_rom[413] = 62;
    assign twf_m0_im_rom[413] = -112;
    assign twf_m0_re_rom[414] = 58;
    assign twf_m0_im_rom[414] = -114;
    assign twf_m0_re_rom[415] = 53;
    assign twf_m0_im_rom[415] = -116;
    assign twf_m0_re_rom[416] = 49;
    assign twf_m0_im_rom[416] = -118;
    assign twf_m0_re_rom[417] = 45;
    assign twf_m0_im_rom[417] = -120;
    assign twf_m0_re_rom[418] = 40;
    assign twf_m0_im_rom[418] = -122;
    assign twf_m0_re_rom[419] = 36;
    assign twf_m0_im_rom[419] = -123;
    assign twf_m0_re_rom[420] = 31;
    assign twf_m0_im_rom[420] = -124;
    assign twf_m0_re_rom[421] = 27;
    assign twf_m0_im_rom[421] = -125;
    assign twf_m0_re_rom[422] = 22;
    assign twf_m0_im_rom[422] = -126;
    assign twf_m0_re_rom[423] = 17;
    assign twf_m0_im_rom[423] = -127;
    assign twf_m0_re_rom[424] = 13;
    assign twf_m0_im_rom[424] = -127;
    assign twf_m0_re_rom[425] = 8;
    assign twf_m0_im_rom[425] = -128;
    assign twf_m0_re_rom[426] = 3;
    assign twf_m0_im_rom[426] = -128;
    assign twf_m0_re_rom[427] = -2;
    assign twf_m0_im_rom[427] = -128;
    assign twf_m0_re_rom[428] = -6;
    assign twf_m0_im_rom[428] = -128;
    assign twf_m0_re_rom[429] = -11;
    assign twf_m0_im_rom[429] = -128;
    assign twf_m0_re_rom[430] = -16;
    assign twf_m0_im_rom[430] = -127;
    assign twf_m0_re_rom[431] = -20;
    assign twf_m0_im_rom[431] = -126;
    assign twf_m0_re_rom[432] = -25;
    assign twf_m0_im_rom[432] = -126;
    assign twf_m0_re_rom[433] = -30;
    assign twf_m0_im_rom[433] = -125;
    assign twf_m0_re_rom[434] = -34;
    assign twf_m0_im_rom[434] = -123;
    assign twf_m0_re_rom[435] = -39;
    assign twf_m0_im_rom[435] = -122;
    assign twf_m0_re_rom[436] = -43;
    assign twf_m0_im_rom[436] = -121;
    assign twf_m0_re_rom[437] = -48;
    assign twf_m0_im_rom[437] = -119;
    assign twf_m0_re_rom[438] = -52;
    assign twf_m0_im_rom[438] = -117;
    assign twf_m0_re_rom[439] = -56;
    assign twf_m0_im_rom[439] = -115;
    assign twf_m0_re_rom[440] = -60;
    assign twf_m0_im_rom[440] = -113;
    assign twf_m0_re_rom[441] = -64;
    assign twf_m0_im_rom[441] = -111;
    assign twf_m0_re_rom[442] = -68;
    assign twf_m0_im_rom[442] = -108;
    assign twf_m0_re_rom[443] = -72;
    assign twf_m0_im_rom[443] = -106;
    assign twf_m0_re_rom[444] = -76;
    assign twf_m0_im_rom[444] = -103;
    assign twf_m0_re_rom[445] = -80;
    assign twf_m0_im_rom[445] = -100;
    assign twf_m0_re_rom[446] = -84;
    assign twf_m0_im_rom[446] = -97;
    assign twf_m0_re_rom[447] = -87;
    assign twf_m0_im_rom[447] = -94;
    assign twf_m0_re_rom[448] = 128;
    assign twf_m0_im_rom[448] = 0;
    assign twf_m0_re_rom[449] = 128;
    assign twf_m0_im_rom[449] = -11;
    assign twf_m0_re_rom[450] = 126;
    assign twf_m0_im_rom[450] = -22;
    assign twf_m0_re_rom[451] = 124;
    assign twf_m0_im_rom[451] = -33;
    assign twf_m0_re_rom[452] = 121;
    assign twf_m0_im_rom[452] = -43;
    assign twf_m0_re_rom[453] = 116;
    assign twf_m0_im_rom[453] = -53;
    assign twf_m0_re_rom[454] = 111;
    assign twf_m0_im_rom[454] = -63;
    assign twf_m0_re_rom[455] = 106;
    assign twf_m0_im_rom[455] = -72;
    assign twf_m0_re_rom[456] = 99;
    assign twf_m0_im_rom[456] = -81;
    assign twf_m0_re_rom[457] = 92;
    assign twf_m0_im_rom[457] = -89;
    assign twf_m0_re_rom[458] = 84;
    assign twf_m0_im_rom[458] = -97;
    assign twf_m0_re_rom[459] = 75;
    assign twf_m0_im_rom[459] = -104;
    assign twf_m0_re_rom[460] = 66;
    assign twf_m0_im_rom[460] = -110;
    assign twf_m0_re_rom[461] = 56;
    assign twf_m0_im_rom[461] = -115;
    assign twf_m0_re_rom[462] = 46;
    assign twf_m0_im_rom[462] = -119;
    assign twf_m0_re_rom[463] = 36;
    assign twf_m0_im_rom[463] = -123;
    assign twf_m0_re_rom[464] = 25;
    assign twf_m0_im_rom[464] = -126;
    assign twf_m0_re_rom[465] = 14;
    assign twf_m0_im_rom[465] = -127;
    assign twf_m0_re_rom[466] = 3;
    assign twf_m0_im_rom[466] = -128;
    assign twf_m0_re_rom[467] = -8;
    assign twf_m0_im_rom[467] = -128;
    assign twf_m0_re_rom[468] = -19;
    assign twf_m0_im_rom[468] = -127;
    assign twf_m0_re_rom[469] = -30;
    assign twf_m0_im_rom[469] = -125;
    assign twf_m0_re_rom[470] = -40;
    assign twf_m0_im_rom[470] = -122;
    assign twf_m0_re_rom[471] = -50;
    assign twf_m0_im_rom[471] = -118;
    assign twf_m0_re_rom[472] = -60;
    assign twf_m0_im_rom[472] = -113;
    assign twf_m0_re_rom[473] = -70;
    assign twf_m0_im_rom[473] = -107;
    assign twf_m0_re_rom[474] = -79;
    assign twf_m0_im_rom[474] = -101;
    assign twf_m0_re_rom[475] = -87;
    assign twf_m0_im_rom[475] = -94;
    assign twf_m0_re_rom[476] = -95;
    assign twf_m0_im_rom[476] = -86;
    assign twf_m0_re_rom[477] = -102;
    assign twf_m0_im_rom[477] = -78;
    assign twf_m0_re_rom[478] = -108;
    assign twf_m0_im_rom[478] = -68;
    assign twf_m0_re_rom[479] = -114;
    assign twf_m0_im_rom[479] = -59;
    assign twf_m0_re_rom[480] = -118;
    assign twf_m0_im_rom[480] = -49;
    assign twf_m0_re_rom[481] = -122;
    assign twf_m0_im_rom[481] = -39;
    assign twf_m0_re_rom[482] = -125;
    assign twf_m0_im_rom[482] = -28;
    assign twf_m0_re_rom[483] = -127;
    assign twf_m0_im_rom[483] = -17;
    assign twf_m0_re_rom[484] = -128;
    assign twf_m0_im_rom[484] = -6;
    assign twf_m0_re_rom[485] = -128;
    assign twf_m0_im_rom[485] = 5;
    assign twf_m0_re_rom[486] = -127;
    assign twf_m0_im_rom[486] = 16;
    assign twf_m0_re_rom[487] = -125;
    assign twf_m0_im_rom[487] = 27;
    assign twf_m0_re_rom[488] = -122;
    assign twf_m0_im_rom[488] = 37;
    assign twf_m0_re_rom[489] = -119;
    assign twf_m0_im_rom[489] = 48;
    assign twf_m0_re_rom[490] = -114;
    assign twf_m0_im_rom[490] = 58;
    assign twf_m0_re_rom[491] = -109;
    assign twf_m0_im_rom[491] = 67;
    assign twf_m0_re_rom[492] = -103;
    assign twf_m0_im_rom[492] = 76;
    assign twf_m0_re_rom[493] = -96;
    assign twf_m0_im_rom[493] = 85;
    assign twf_m0_re_rom[494] = -88;
    assign twf_m0_im_rom[494] = 93;
    assign twf_m0_re_rom[495] = -80;
    assign twf_m0_im_rom[495] = 100;
    assign twf_m0_re_rom[496] = -71;
    assign twf_m0_im_rom[496] = 106;
    assign twf_m0_re_rom[497] = -62;
    assign twf_m0_im_rom[497] = 112;
    assign twf_m0_re_rom[498] = -52;
    assign twf_m0_im_rom[498] = 117;
    assign twf_m0_re_rom[499] = -42;
    assign twf_m0_im_rom[499] = 121;
    assign twf_m0_re_rom[500] = -31;
    assign twf_m0_im_rom[500] = 124;
    assign twf_m0_re_rom[501] = -20;
    assign twf_m0_im_rom[501] = 126;
    assign twf_m0_re_rom[502] = -9;
    assign twf_m0_im_rom[502] = 128;
    assign twf_m0_re_rom[503] = 2;
    assign twf_m0_im_rom[503] = 128;
    assign twf_m0_re_rom[504] = 13;
    assign twf_m0_im_rom[504] = 127;
    assign twf_m0_re_rom[505] = 23;
    assign twf_m0_im_rom[505] = 126;
    assign twf_m0_re_rom[506] = 34;
    assign twf_m0_im_rom[506] = 123;
    assign twf_m0_re_rom[507] = 45;
    assign twf_m0_im_rom[507] = 120;
    assign twf_m0_re_rom[508] = 55;
    assign twf_m0_im_rom[508] = 116;
    assign twf_m0_re_rom[509] = 64;
    assign twf_m0_im_rom[509] = 111;
    assign twf_m0_re_rom[510] = 74;
    assign twf_m0_im_rom[510] = 105;
    assign twf_m0_re_rom[511] = 82;
    assign twf_m0_im_rom[511] = 98;

endmodule
